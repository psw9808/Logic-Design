module findD(input[6:0] p,q,input[13:0] e, output reg[13:0] d);
	integer i,phi;
	
	always@(*) begin
	phi = (p-1)*(q-1);
		if((e*2)%phi==1) d = 2;
		else if((e*3)%phi==1) d = 3;
		else if((e*5)%phi==1) d = 5;
		else if((e*7)%phi==1) d = 7;
		else if((e*11)%phi==1) d = 11;
		else if((e*13)%phi==1) d = 13;
		else if((e*17)%phi==1) d = 17;
		else if((e*19)%phi==1) d = 19;
		else if((e*23)%phi==1) d = 23;
		else if((e*29)%phi==1) d = 29;
		else if((e*31)%phi==1) d = 31;
		else if((e*37)%phi==1) d = 37;
		else if((e*41)%phi==1) d = 41;
		else if((e*43)%phi==1) d = 43;
		else if((e*47)%phi==1) d = 47;
		else if((e*53)%phi==1) d = 53;
		else if((e*59)%phi==1) d = 59;
		else if((e*61)%phi==1) d = 61;
		else if((e*67)%phi==1) d = 67;
		else if((e*71)%phi==1) d = 71;
		else if((e*73)%phi==1) d = 73;
		else if((e*79)%phi==1) d = 79;
		else if((e*83)%phi==1) d = 83;
		else if((e*89)%phi==1) d = 89;
		else if((e*97)%phi==1) d = 97;
		else if((e*101)%phi==1) d = 101;
		else if((e*103)%phi==1) d = 103;
		else if((e*107)%phi==1) d = 107;
		else if((e*109)%phi==1) d = 109;
		else if((e*113)%phi==1) d = 113;
		else if((e*127)%phi==1) d = 127;
		else if((e*131)%phi==1) d = 131;
		else if((e*137)%phi==1) d = 137;
		else if((e*139)%phi==1) d = 139;
		else if((e*149)%phi==1) d = 149;
		else if((e*151)%phi==1) d = 151;
		else if((e*157)%phi==1) d = 157;
		else if((e*163)%phi==1) d = 163;
		else if((e*167)%phi==1) d = 167;
		else if((e*173)%phi==1) d = 173;
		else if((e*179)%phi==1) d = 179;
		else if((e*181)%phi==1) d = 181;
		else if((e*191)%phi==1) d = 191;
		else if((e*193)%phi==1) d = 193;
		else if((e*197)%phi==1) d = 197;
		else if((e*199)%phi==1) d = 199;
		else if((e*211)%phi==1) d = 211;
		else if((e*223)%phi==1) d = 223;
		else if((e*227)%phi==1) d = 227;
		else if((e*229)%phi==1) d = 229;
		else if((e*233)%phi==1) d = 233;
		else if((e*239)%phi==1) d = 239;
		else if((e*241)%phi==1) d = 241;
		else if((e*251)%phi==1) d = 251;
		else if((e*257)%phi==1) d = 257;
		else if((e*263)%phi==1) d = 263;
		else if((e*269)%phi==1) d = 269;
		else if((e*271)%phi==1) d = 271;
		else if((e*277)%phi==1) d = 277;
		else if((e*281)%phi==1) d = 281;
		else if((e*283)%phi==1) d = 283;
		else if((e*293)%phi==1) d = 293;
		else if((e*307)%phi==1) d = 307;
		else if((e*311)%phi==1) d = 311;
		else if((e*313)%phi==1) d = 313;
		else if((e*317)%phi==1) d = 317;
		else if((e*331)%phi==1) d = 331;
		else if((e*337)%phi==1) d = 337;
		else if((e*347)%phi==1) d = 347;
		else if((e*349)%phi==1) d = 349;
		else if((e*353)%phi==1) d = 353;
		else if((e*359)%phi==1) d = 359;
		else if((e*367)%phi==1) d = 367;
		else if((e*373)%phi==1) d = 373;
		else if((e*379)%phi==1) d = 379;
		else if((e*383)%phi==1) d = 383;
		else if((e*389)%phi==1) d = 389;
		else if((e*397)%phi==1) d = 397;
		else if((e*401)%phi==1) d = 401;
		else if((e*409)%phi==1) d = 409;
		else if((e*419)%phi==1) d = 419;
		else if((e*421)%phi==1) d = 421;
		else if((e*431)%phi==1) d = 431;
		else if((e*433)%phi==1) d = 433;
		else if((e*439)%phi==1) d = 439;
		else if((e*443)%phi==1) d = 443;
		else if((e*449)%phi==1) d = 449;
		else if((e*457)%phi==1) d = 457;
		else if((e*461)%phi==1) d = 461;
		else if((e*463)%phi==1) d = 463;
		else if((e*467)%phi==1) d = 467;
		else if((e*479)%phi==1) d = 479;
		else if((e*487)%phi==1) d = 487;
		else if((e*491)%phi==1) d = 491;
		else if((e*499)%phi==1) d = 499;
		else if((e*503)%phi==1) d = 503;
		else if((e*509)%phi==1) d = 509;
		else if((e*521)%phi==1) d = 521;
		else if((e*523)%phi==1) d = 523;
		else if((e*541)%phi==1) d = 541;
		else if((e*547)%phi==1) d = 547;
		else if((e*557)%phi==1) d = 557;
		else if((e*563)%phi==1) d = 563;
		else if((e*569)%phi==1) d = 569;
		else if((e*571)%phi==1) d = 571;
		else if((e*577)%phi==1) d = 577;
		else if((e*587)%phi==1) d = 587;
		else if((e*593)%phi==1) d = 593;
		else if((e*599)%phi==1) d = 599;
		else if((e*601)%phi==1) d = 601;
		else if((e*607)%phi==1) d = 607;
		else if((e*613)%phi==1) d = 613;
		else if((e*617)%phi==1) d = 617;
		else if((e*619)%phi==1) d = 619;
		else if((e*631)%phi==1) d = 631;
		else if((e*641)%phi==1) d = 641;
		else if((e*643)%phi==1) d = 643;
		else if((e*647)%phi==1) d = 647;
		else if((e*653)%phi==1) d = 653;
		else if((e*659)%phi==1) d = 659;
		else if((e*661)%phi==1) d = 661;
		else if((e*673)%phi==1) d = 673;
		else if((e*677)%phi==1) d = 677;
		else if((e*683)%phi==1) d = 683;
		else if((e*691)%phi==1) d = 691;
		else if((e*701)%phi==1) d = 701;
		else if((e*709)%phi==1) d = 709;
		else if((e*719)%phi==1) d = 719;
		else if((e*727)%phi==1) d = 727;
		else if((e*733)%phi==1) d = 733;
		else if((e*739)%phi==1) d = 739;
		else if((e*743)%phi==1) d = 743;
		else if((e*751)%phi==1) d = 751;
		else if((e*757)%phi==1) d = 757;
		else if((e*761)%phi==1) d = 761;
		else if((e*769)%phi==1) d = 769;
		else if((e*773)%phi==1) d = 773;
		else if((e*787)%phi==1) d = 787;
		else if((e*797)%phi==1) d = 797;
		else if((e*809)%phi==1) d = 809;
		else if((e*811)%phi==1) d = 811;
		else if((e*821)%phi==1) d = 821;
		else if((e*823)%phi==1) d = 823;
		else if((e*827)%phi==1) d = 827;
		else if((e*829)%phi==1) d = 829;
		else if((e*839)%phi==1) d = 839;
		else if((e*853)%phi==1) d = 853;
		else if((e*857)%phi==1) d = 857;
		else if((e*859)%phi==1) d = 859;
		else if((e*863)%phi==1) d = 863;
		else if((e*877)%phi==1) d = 877;
		else if((e*881)%phi==1) d = 881;
		else if((e*883)%phi==1) d = 883;
		else if((e*887)%phi==1) d = 887;
		else if((e*907)%phi==1) d = 907;
		else if((e*911)%phi==1) d = 911;
		else if((e*919)%phi==1) d = 919;
		else if((e*929)%phi==1) d = 929;
		else if((e*937)%phi==1) d = 937;
		else if((e*941)%phi==1) d = 941;
		else if((e*947)%phi==1) d = 947;
		else if((e*953)%phi==1) d = 953;
		else if((e*967)%phi==1) d = 967;
		else if((e*971)%phi==1) d = 971;
		else if((e*977)%phi==1) d = 977;
		else if((e*983)%phi==1) d = 983;
		else if((e*991)%phi==1) d = 991;
		else if((e*997)%phi==1) d = 997;
		else if((e*1009)%phi==1) d = 1009;
		else if((e*1013)%phi==1) d = 1013;
		else if((e*1019)%phi==1) d = 1019;
		else if((e*1021)%phi==1) d = 1021;
		else if((e*1031)%phi==1) d = 1031;
		else if((e*1033)%phi==1) d = 1033;
		else if((e*1039)%phi==1) d = 1039;
		else if((e*1049)%phi==1) d = 1049;
		else if((e*1051)%phi==1) d = 1051;
		else if((e*1061)%phi==1) d = 1061;
		else if((e*1063)%phi==1) d = 1063;
		else if((e*1069)%phi==1) d = 1069;
		else if((e*1087)%phi==1) d = 1087;
		else if((e*1091)%phi==1) d = 1091;
		else if((e*1093)%phi==1) d = 1093;
		else if((e*1097)%phi==1) d = 1097;
		else if((e*1103)%phi==1) d = 1103;
		else if((e*1109)%phi==1) d = 1109;
		else if((e*1117)%phi==1) d = 1117;
		else if((e*1123)%phi==1) d = 1123;
		else if((e*1129)%phi==1) d = 1129;
		else if((e*1151)%phi==1) d = 1151;
		else if((e*1153)%phi==1) d = 1153;
		else if((e*1163)%phi==1) d = 1163;
		else if((e*1171)%phi==1) d = 1171;
		else if((e*1181)%phi==1) d = 1181;
		else if((e*1187)%phi==1) d = 1187;
		else if((e*1193)%phi==1) d = 1193;
		else if((e*1201)%phi==1) d = 1201;
		else if((e*1213)%phi==1) d = 1213;
		else if((e*1217)%phi==1) d = 1217;
		else if((e*1223)%phi==1) d = 1223;
		
		else begin
			for(i=4095; i>1224; i=i-2) begin
				if((e*i)%phi==1)begin
					d = i;
				end
			end
		end
		
	end
endmodule