module sub(output[15:0] z, input[15:0] a,b);
	assign z=a-b;
endmodule
