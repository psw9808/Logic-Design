module mul(input[15:0] a,b, output[15:0] out, output overflow);
	wire[15:0] a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15;
	wire[15:0] o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14;
	wire c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15;
	wire r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r16,r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28;
	
	multiandgate u0(a,b[0],a0);
	multiandgate u1(a,b[1],a1);
	multiandgate u2(a,b[2],a2);
	multiandgate u3(a,b[3],a3);
	multiandgate u4(a,b[4],a4);
	multiandgate u5(a,b[5],a5);
	multiandgate u6(a,b[6],a6);
	multiandgate u7(a,b[7],a7);
	multiandgate u8(a,b[8],a8);
	multiandgate u9(a,b[9],a9);
	multiandgate u10(a,b[10],a10);
	multiandgate u11(a,b[11],a11);
	multiandgate u12(a,b[12],a12);
	multiandgate u13(a,b[13],a13);
	multiandgate u14(a,b[14],a14);
	multiandgate u15(a,b[15],a15);
	
	bit16adder add0(a0, a1<<1, 0, o1, c1);
	bit16adder add1(o1, a2<<2, 0, o2, c2);
	bit16adder add2(o2, a3<<3, 0, o3, c3);
	bit16adder add3(o3, a4<<4, 0, o4, c4);
	bit16adder add4(o4, a5<<5, 0, o5, c5);
	bit16adder add5(o5, a6<<6, 0, o6, c6);
	bit16adder add6(o6, a7<<7, 0, o7, c7);
	bit16adder add7(o7, a8<<8, 0, o8, c8);
	bit16adder add8(o8, a9<<9, 0, o9, c9);
	bit16adder add9(o9, a10<<10, 0, o10, c10);
	bit16adder add10(o10, a11<<11, 0, o11, c11);
	bit16adder add11(o11, a12<<12, 0, o12, c12);
	bit16adder add12(o12, a13<<13, 0, o13, c13);
	bit16adder add13(o13, a14<<14, 0, o14, c14);
	bit16adder add14(o14, a15<<15, 0, out, c15);
	
	or or1(r1,|(a15>>1),|(a14>>2));
	or or2(r2,r1,|(a13>>3));
	or or3(r3,r2,|(a12>>4));
	or or4(r4,r3,|(a11>>5));
	or or5(r5,r4,|(a10>>6));
	or or6(r6,r5,|(a9>>7));
	or or7(r7,r6,|(a8>>8));
	or or8(r8,r7,|(a7>>9));
	or or9(r9,r8,|(a6>>10));
	or or10(r10,r9,|(a5>>11));
	or or11(r11,r10,|(a4>>12));
	or or12(r12,r11,|(a3>>13));
	or or13(r13,r12,|(a2>>14));
	or or14(r14,r13,|(a1>>15));
	or or15(r15,r14,c1);
	or or16(r16,r15,c2);
	or or17(r17,r16,c3);
	or or18(r18,r17,c4);
	or or19(r19,r18,c5);
	or or20(r20,r19,c6);
	or or21(r21,r20,c7);
	or or22(r22,r21,c8);
	or or23(r23,r22,c9);
	or or24(r24,r23,c10);
	or or25(r25,r24,c11);
	or or26(r26,r25,c12);
	or or27(r27,r26,c13);
	or or28(r28,r27,c14);
	or or29(overflow,r28,c15);
	
endmodule